
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Ram1 is
    Port ( 
				clock 	: in  	std_logic;
		--		reset 	: in  	std_logic;
				address1 	: in 		std_logic_vector(11 downto 0);
				data1 	: out 	std_logic_vector(3 downto 0)

		
			  );
end Ram1;

architecture Behavioral of Ram1 is

component RAMB16_S4_S4 is
generic( 	INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
				);
port(
		WEA  : in std_logic;
		ENA  : in std_logic;
		SSRA : in std_logic;
		CLKA : in std_logic;
		ADDRA: in std_logic_vector(11 downto 0);
		DIA  : in std_logic_vector(3 downto 0);
		DOA  : out std_logic_vector(3 downto 0);
		
		WEB  : in std_logic;
		ENB  : in std_logic;
		SSRB : in std_logic;
		CLKB : in std_logic;
		ADDRB: in std_logic_vector(11 downto 0);
		DIB  : in std_logic_vector(3 downto 0);
		DOB  : out std_logic_vector(3 downto 0)
		);
end component;

signal dummy : std_logic_vector( 3 downto 0);

	begin
		MEM: RAMB16_S4_S4
		generic map(

		--Marlin1  0~2431
      INIT_00 => X"8888888888888888888888886646664565888888888888888888888888888888",
      INIT_01 => X"8888888888888888888888866644044555888888888888888888888888888888",
      INIT_02 => X"8888888888888888888888666001111105588888888888888888888888888888",
      INIT_03 => X"8888888888888888888845111111111115588888888888888888888888888888",
      INIT_04 => X"8888888888888888888811111111111140588888888888888888888888888888",
      INIT_05 => X"8888888888888888861111111111111111058888888888888888888888888888",
      INIT_06 => X"8888888888888888845111111111111111558888888888888888888888888888",
      INIT_07 => X"8888888888888886451111111111111111057888888888888888888888888888",
      INIT_08 => X"8888888888888846661111111111111111058888888888888888888888888888",
      INIT_09 => X"8888888888884677761111111111111111158888888888888888888888888888",
      INIT_0A => X"8888888888846556000611111111111115555888888888888888888888888888",
      INIT_0B => X"8888888884511111566651111111111146655668888888888888888888888888",
      INIT_0C => X"8888886451111111156665111111111166665555555888888888888888888888",
      INIT_0D => X"8888866611111111111566511111111106661111155558888888888888888888",
      INIT_0E => X"8888885111111111111166651111111104666111111145555888888888888888",
      INIT_0F => X"8888855111111111111114665111111016666011111115555888888888888888",
      INIT_10 => X"8884455111111111111110665111110466666001111111155888888888888888",
      INIT_11 => X"8887650111155511111110665111110466666605511111155888888888888888",
      INIT_12 => X"6888656111007751111111466111104666666605555111114588888888644448",
      INIT_13 => X"8888661115007775111111466111114666666660555551156688888644805118",
      INIT_14 => X"8888611116567775111111566111166666666655555551156888800055111118",
		INIT_15 => X"8885111177777665111111566514666666666655555555660008511111111118",
      INIT_16 => X"8885111115777775111110664114666666666505555566666511111111111118",
      INIT_17 => X"8885111111577751111111146411166666665115055566666611111111111118",
      INIT_18 => X"8881111111111111111115516411166666451111505556666641111111111448",
      INIT_19 => X"8881111111111111111111146411166665511111150554666641111111111488",
      INIT_1A => X"8881111111111111111111146411104111111111115055466611111111111488",
		INIT_1B => X"8886111111111111111111156411111111111111110554666115151511111488",
      INIT_1C => X"8885100001111111111111156451111111111111111055466665155555111488",
      INIT_1D => X"8885110000005111111111556145511111111111111115546666555555111488",
      INIT_1E => X"8888511111111111111111146555551111111111111105546666055555111488",
      INIT_1F => X"8888811111151515151515546551515111111111111050546646455555111118",
      INIT_20 => X"8888881111515151115151155465050551111111115055056666451555511118",
      INIT_21 => X"8888885111151115111155566555555551111111115050546666455151111111",
      INIT_22 => X"8888888886655665566666665555515151111111150550541644445151111118",
      INIT_23 => X"8888888888846586665651151554551555111111505050504440048848841118",
      INIT_24 => X"8888888888888885151515151151515156111115150505044488848884888844",
      INIT_25 => X"8888888888888888888855555488851515155558856888888888888888888888",
		
		--heart 2432~2879
--		88881118888881118888
--		88811111188111111888
--		88111111188111111188
--		81111111111111111118
--		81111111111111111118
--		11111111111111111111
--		11111111111111111111
--		11111111111111111111
--		11111111111111111111
--		81111111111111111118
--		81111111111111111118
--		88111111111111111188
--		88111111111111111188
--		88811111111111111888
--		88811111111111111888
--		88881111111111118888
--		88888111111111188888
--		88888881111111888888
--		88888888811888888888
--		88888888888888888888
		INIT_26 => X"8888111888888111888888811111188111111888881111111881111111888111",
		INIT_27 => X"1111111111111118811111111111111111181111111111111111111111111111",
		INIT_28 => X"1111111111111111111111111111111111111111111111111111811111111111",
		INIT_29 => X"1111111881111111111111111118881111111111111111888811111111111111",
		INIT_2A => X"1188888111111111111118888881111111111111188888881111111111118888",
		INIT_2B => X"8888811111111118888888888881111111888888888888888118888888888888",
		INIT_2C => X"8888888888888888000000000000000000000000000000000000000000000000",		
		--! 2880~3327
--		88888880000008888888
--		88880333333333308888
--		88033333333333333088
--		03333333333333333330
--		03333333333333333330
--		80333333333333333308
--		80333333333333333308
--		80333333333333333308
--		80333333333333333308
--		88033333333333333088
--		88803333333333330888
--		88880333333333008888
--		88888033333333088888
--		88888880000008888888
--		88888888888888888888
--		88888888800888888888
--		88888888033088888888
--		88888888033088888888
--		88888888800888888888
--		88888888888888888888

		INIT_2D => X"8888888000000888888888880333333333308888880333333333333330880333",
		INIT_2E => X"3333333333333330033333333333333333308033333333333333330880333333",
		INIT_2F => X"3333333333088033333333333333330880333333333333333308880333333333",
		INIT_30 => X"3333308888803333333333330888888803333333330088888888803333333308",
		INIT_31 => X"8888888888800000088888888888888888888888888888888888800888888888",
		INIT_32 => X"8888888803308888888888888888033088888888888888888008888888888888",
		INIT_33 => X"8888888888888888000000000000000000000000000000000000000000000000",
      
    
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
						WEA => '0',				-- I never need to write to A, just read from it
						ENA  => '1',			-- Always enable A for reading
						SSRA => '0',			-- set to 0
						CLKA => clock,			-- take the clock coming from the top level
						ADDRA => address1,			-- address comes in from rgb_reader
						DIA  => "0111",
						DOA  => data1, 
						
						WEB => '0',				
						ENB  => '0',
						SSRB => '0',
						CLKB => clock,
						ADDRB => "000000000000",
						DIB  => "0111",
						DOB  => dummy
				);					
				
end Behavioral;
