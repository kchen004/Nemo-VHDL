
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Ram2 is
    Port ( 
				clock 	: in  	std_logic;
				address 	: in 		std_logic_vector(11 downto 0);
				data  	: out  	std_logic_vector(3 downto 0)
		
			  );
end Ram2;

architecture Behavioral of Ram2 is

component RAMB16_S4_S4 is
generic( 	INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
				);
port(
		WEA  : in std_logic;
		ENA  : in std_logic;
		SSRA : in std_logic;
		CLKA : in std_logic;
		ADDRA: in std_logic_vector(11 downto 0);
		DIA  : in std_logic_vector(3 downto 0);
		DOA  : out std_logic_vector(3 downto 0);
		
		WEB  : in std_logic;
		ENB  : in std_logic;
		SSRB : in std_logic;
		CLKB : in std_logic;
		ADDRB: in std_logic_vector(11 downto 0);
		DIB  : in std_logic_vector(3 downto 0);
		DOB  : out std_logic_vector(3 downto 0)
		);
end component;

signal dummy : std_logic_vector( 3 downto 0);

	begin
		MEM: RAMB16_S4_S4
		generic map(
		
		--Jellyfish
	
		INIT_00 => X"8888888888888888888888888000088888888888888888888888888888888888",
      INIT_01 => X"8888888888888888888888460000440060888888888888888888888888888888",
      INIT_02 => X"8888888888888888804604604060460460460460406488888888888888888888",
      INIT_03 => X"8888888888888888804604604060460460460460406488888888888888888888",
      INIT_04 => X"8888888888888804604464646464646464644640406404688888888888888888",
      INIT_05 => X"8888888888888804604464646464646464644640406404688888888888888888",
      INIT_06 => X"8888888888804604646464646464646464646464646404608888888888888888",
      INIT_07 => X"8888888888804604446146166616661666166441646446608888888888888888",
      INIT_08 => X"8888888804046044461461666166616661664416464466408888888888888888",
      INIT_09 => X"8888884004046044461461666166666661664416464466408888888888888888",
      INIT_0A => X"8888884004046044461461666666616661664416464466408888888888888888",
      INIT_0B => X"8880404004046044461461666666316661663416464466408888888888888888",
      INIT_0C => X"8880404004046044461461366666316661663416464466408888888888888888",
      INIT_0D => X"8804404004046044461461663336316661663416464666408888888888888888",
      INIT_0E => X"8043600084446660003656056056056600606003400000888888888888888888",
      INIT_0F => X"0044448563565654661565656565655444063464360080888888888888888888",
      INIT_10 => X"0003636363463636361366346436366366435834630088888888888888888888",
      INIT_11 => X"0000000000000000000444444000000000000000888888888888888888888888",
      INIT_12 => X"8800000000000000000000000000000000000008888888888888888888888888",
      INIT_13 => X"8880000000000000000000000000000000000888888888888888888888888888",
      INIT_14 => X"8888000000000000000000000000000000888888888888888888888888888888",
      INIT_15 => X"8888888888887778878877888888888777888888888888888888888888888888",
      INIT_16 => X"8888888888887778877887788888887778888888888888888888888888888888",
      INIT_17 => X"8888888888887778778880788888878778888888888888888888888888888888",
      INIT_18 => X"8888888888877888788888708888807888888888888888888888888888888888",
      INIT_19 => X"8888888888877887888888778888778888888888888888888888888888888888",
      INIT_1A => X"8888888888777887888887078880708888888888888888888888888888888888",
      INIT_1B => X"8888888877078807888870770788807888888888888888888888888888888888",
      INIT_1C => X"8888888707888880788778888888887078888888888888888888888888888888",
      INIT_1D => X"8888877788888878700788888888870788888888888888888888888888888888",
      INIT_1E => X"8888778888888878870888888888788888888888888888888888888888888888",
		INIT_1F => X"8887088888887878807888888888088888888888888888888888888888888888",
      INIT_20 => X"7778888888887888880788888888807888888888888888888888888888888888",
      INIT_21 => X"8888888888887888888877888888708888888888888888888888888888888888",
      INIT_22 => X"8888888888887888888887888888877888888888888888888888888888888888",
      INIT_23 => X"8888888888887888888887788888880888888888888888888888888888888888",
      INIT_24 => X"8888888888870888888778888888887788888888888888888888888888888888",
		INIT_25 => X"8888888888870888887888888888878888888888888888888888888888888888",
      INIT_26 => X"8888888880788888878888888888870888888888888888888888888888888888",
      INIT_27 => X"8888888700888878788788888888708888888888888888888888888888888888",
      INIT_28 => X"8888887778888888888888888888708888888888888888888888888888888888",
      INIT_29 => X"8888877888888888888888888880788888888888888888888888888888888888",
      INIT_2A => X"8888788888888888888888888888778888888888888888888888888888888888",
      INIT_2B => X"8888788888888888888888888777788888888888888888888888888888888888",
      INIT_2C => X"8888777888888888888888887788888888888888888888888888888888888888",
      INIT_2D => X"8888888888888888888888078888888888888888888888888888888888888888",
      INIT_2E => X"8888888888888888888887088888888888888888888888888888888888888888",
      INIT_2F => X"8888888888888888888887888888888888888888888888888888888888888888",
      INIT_30 => X"8888888888888888887788888888888888888888888888888888888888888888",
      INIT_31 => X"8888888888888888878888888888888888888888888888888888888888888888",
		
		
		
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      
		
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
						WEA => '0',				-- I never need to write to A, just read from it
						ENA  => '1',			-- Always enable A for reading
						SSRA => '0',			-- set to 0
						CLKA => clock,			-- take the clock coming from the top level
						ADDRA => address,			-- address comes in from rgb_reader
						DIA  => "0111",
						DOA  => data, 
						
						WEB => '0',				
						ENB  => '0',
						SSRB => '0',
						CLKB => clock,
						ADDRB => "000000000000",
						DIB  =>  "0000",
						DOB  => dummy
				);					
				
end Behavioral;
