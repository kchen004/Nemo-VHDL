library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity enemy_ram is
    Port ( 
				clk 	: in  	std_logic;

				portA_address 	: in 		std_logic_vector(8 downto 0);
				portA_dataIn  	: in  	std_logic_vector(31 downto 0);
				portA_dataOut  : out 	std_logic_vector(31 downto 0);
				portA_write		: in		std_logic;
				
				portB_address 	: in 		std_logic_vector(8 downto 0);
				portB_data  	: out  	std_logic_vector(31 downto 0)
		
			  );
end enemy_ram;

   -- RAMB16_S36_S36: Virtex-II/II-Pro, Spartan-3/3E 512 x 32 + 4 Parity bits Dual-Port RAM
   -- Xilinx HDL Language Template, version 9.1i

architecture Behavioral of enemy_ram is

component   RAMB16_S36_S36 is
   generic(	INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
				INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000");
   port (
      DOA 	: out std_logic_vector (31 downto 0);      -- Port A 32-bit Data Output
      DOB 	: out std_logic_vector (31 downto 0);      -- Port B 32-bit Data Output
      DOPA 	: out std_logic_vector (3 downto 0);     -- Port A 4-bit Parity Output
      DOPB 	: out std_logic_vector (3 downto 0);     -- Port B 4-bit Parity Output
      ADDRA : in std_logic_vector (8 downto 0);   -- Port A 9-bit Address Input
      ADDRB : in std_logic_vector (8 downto 0);   -- Port B 9-bit Address Input
      CLKA 	: in std_logic;    -- Port A Clock
      CLKB 	: in std_logic;    -- Port B Clock
      DIA 	: in std_logic_vector (31 downto 0);        -- Port A 32-bit Data Input
      DIB 	: in std_logic_vector (31 downto 0);        -- Port B 32-bit Data Input
      DIPA 	: in std_logic_vector (3 downto 0);    -- Port A 4-bit parity Input
      DIPB 	: in std_logic_vector (3 downto 0);    -- Port-B 4-bit parity Input
      ENA  	: in std_logic;      -- Port A RAM Enable Input
      ENB 	: in std_logic;      -- PortB RAM Enable Input
      SSRA 	: in std_logic;    -- Port A Synchronous Set/Reset Input
      SSRB 	: in std_logic;    -- Port B Synchronous Set/Reset Input
      WEA 	: in std_logic;     -- Port A Write Enable Input
      WEB 	: in std_logic  -- Port B Write Enable Input
   );

   -- End of RAMB16_S36_S36_inst instantiation
end component;

signal dummy1 : std_logic_vector( 3 downto 0);
signal dummy2 : std_logic_vector( 3 downto 0);

	begin
		E_MEM: RAMB16_S36_S36
	--	generic map(
	--	)

				port map (
					DOA => portA_dataOut,      -- Port A 32-bit Data Output
					DOB => portB_data,      -- Port B 32-bit Data Output
					DOPA => dummy1,    -- Port A 4-bit Parity Output
					DOPB => dummy2,    -- Port B 4-bit Parity Output
					ADDRA => portA_address,  -- Port A 9-bit Address Input
					ADDRB => portB_address,  -- Port B 9-bit Address Input
					CLKA => clk,    -- Port A Clock
					CLKB => clk,    -- Port B Clock
					DIA => portA_dataIn,      -- Port A 32-bit Data Input
					DIB => "00000000000000000000000000000000",      -- Port B 32-bit Data Input
					DIPA => "0000",    -- Port A 4-bit parity Input
					DIPB => "0000",    -- Port-B 4-bit parity Input
					ENA => '1',      -- Port A RAM Enable Input
					ENB => '1',      -- PortB RAM Enable Input
					SSRA => '0',    -- Port A Synchronous Set/Reset Input
					SSRB => '0',    -- Port B Synchronous Set/Reset Input
					WEA => portA_write,      -- Port A Write Enable Input
					WEB => '0'       -- Port B Write Enable Input
				);					
				
end Behavioral;

